/*
 *
 *
 *
 *
 *
 *
 */
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.types.all;
use work.all;


entity test_bench is
end test_bench;


architecture test of test_bench is



begin

    

end test;
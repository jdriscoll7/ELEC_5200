/* File: register.v
 * 
 * Implements a generic register model.
 *
 */
 

module register #(parameter SIZE = 8) 
                 (input  [(SIZE-1):0] data_in,
                  output [(SIZE-1):0] data_out
                  input               clock);

endmodule

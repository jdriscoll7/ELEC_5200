/* File: control_unit.v
 *
 * - Implements the controller used in the CPU design. Essentially
 *   coordinates all of the control signals for datapath.
 *
 */


/* Module for the control unit.
 *  
 * - Inputs:
 *     - op_code: 4 bit opcode from instruction 
 *
 *
 *
 *
 *
 */
module control_unit (input [3:0] op_code,
                     input [1:0] cond);
 
 
 
endmodule
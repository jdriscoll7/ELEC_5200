/* File: control_unit.v
 *
 * - Implements the controller used in the CPU design. Essentially
 *   coordinates all of the control signals for datapath.
 *
 */


/* Module for the control unit.
 *  
 * - Inputs:
 *     - op_code: 4-bit opcode from instruction
 *     - cond:    2-bit conditional code from branch instructions
 *
 * - Outputs:
 *     - 
 *
 *
 *
 *
 */
module control_unit (input [3:0] op_code,
                     input [1:0] cond);
 
 
 
endmodule